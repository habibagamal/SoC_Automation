module ana (PAD);
    inout PAD;
endmodule