module do (out, PAD);
    input out;
    output PAD;

    assign PAD = out;
endmodule